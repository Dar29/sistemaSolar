--------------------------------------------------------------------------------
-- Nombre: Jose Diaz
-- Fecha:  9/10/2024
--------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity Compuerta1 is
    Port (	e1: in STD_LOGIC;
			e2: in STD_LOGIC;
			s:  out STD_LOGIC; 	            
);
end Compuerta1 ;

architecture Behavioral of Compuerta1 is
– COMPONENTS
– SIGNALS

begin
– DISEÑO

end Behavioral;
