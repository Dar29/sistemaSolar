--------------------------------------------------------------------------------
-- Nombre: Nombre del creador
-- Fecha:  dia/mes/año
--------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity <Entidad> is
    Port (	<entrada1>: in STD_LOGIC;
			<entrada2>: in STD_LOGIC_VECTOR (7 downto 0);
			<salida1>:  out STD_LOGIC; 	
			<salida2>:  out STD_LOGIC_VECTOR (7 downto 0)              
);
end <Entidad> ;

architecture Behavioral of <Entidad>  is
-- COMPONENTS
-- SIGNALS

begin
-- DISEÑO

end Behavioral;
